module ctrl(
    output reg_write, 
    output [3:0] aluop, 
    input [5:0] op, 
    input funct);

endmodule
